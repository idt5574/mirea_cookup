         42 merch�            kyrit_kruto�.           Goblin@B          Wok�            Burger�       